magic
tech sky130A
magscale 1 2
timestamp 1717266104
<< metal1 >>
rect 19667 11650 19673 11702
rect 19725 11694 19731 11702
rect 19725 11658 19767 11694
rect 19725 11650 19731 11658
rect 29695 11546 29701 11554
rect 29659 11510 29701 11546
rect 29695 11502 29701 11510
rect 29753 11502 29759 11554
rect 29695 11176 29701 11184
rect 29659 11140 29701 11176
rect 29695 11132 29701 11140
rect 29753 11132 29759 11184
rect 19567 10910 19573 10962
rect 19625 10954 19631 10962
rect 19625 10918 19767 10954
rect 19625 10910 19631 10918
rect 19667 10392 19673 10444
rect 19725 10436 19731 10444
rect 19725 10400 19767 10436
rect 19725 10392 19731 10400
rect 29695 10214 29701 10222
rect 29659 10178 29701 10214
rect 29695 10170 29701 10178
rect 29753 10170 29759 10222
rect 29695 9844 29701 9852
rect 29659 9808 29701 9844
rect 29695 9800 29701 9808
rect 29753 9800 29759 9852
rect 19567 9578 19573 9630
rect 19625 9622 19631 9630
rect 19625 9586 19767 9622
rect 19625 9578 19631 9586
rect 19667 9060 19673 9112
rect 19725 9104 19731 9112
rect 19725 9068 19767 9104
rect 19725 9060 19731 9068
rect 29695 8882 29701 8890
rect 29659 8846 29701 8882
rect 29695 8838 29701 8846
rect 29753 8838 29759 8890
rect 29695 8512 29701 8520
rect 29659 8476 29701 8512
rect 29695 8468 29701 8476
rect 29753 8468 29759 8520
rect 19567 8246 19573 8298
rect 19625 8290 19631 8298
rect 19625 8254 19767 8290
rect 19625 8246 19631 8254
rect 19667 7728 19673 7780
rect 19725 7772 19731 7780
rect 19725 7736 19767 7772
rect 19725 7728 19731 7736
rect 29695 7550 29701 7558
rect 29659 7514 29701 7550
rect 29695 7506 29701 7514
rect 29753 7506 29759 7558
rect 29695 7180 29701 7188
rect 29659 7144 29701 7180
rect 29695 7136 29701 7144
rect 29753 7136 29759 7188
rect 19567 6914 19573 6966
rect 19625 6958 19631 6966
rect 19625 6922 19767 6958
rect 19625 6914 19631 6922
rect 13678 4034 13684 4035
rect 13361 3984 13684 4034
rect 13678 3983 13684 3984
rect 13736 3983 13742 4035
rect 20254 1960 20306 2000
rect 20358 1960 20410 2000
rect 29086 1960 29138 2000
rect 29190 1960 29242 2000
rect 19994 1840 20254 1960
rect 20306 1840 20312 1960
rect 20352 1840 20358 1960
rect 20410 1840 20670 1960
rect 28826 1840 29086 1960
rect 29138 1840 29144 1960
rect 29184 1840 29190 1960
rect 29242 1840 29502 1960
<< via1 >>
rect 19673 11650 19725 11702
rect 29701 11502 29753 11554
rect 29701 11132 29753 11184
rect 19573 10910 19625 10962
rect 19673 10392 19725 10444
rect 29701 10170 29753 10222
rect 29701 9800 29753 9852
rect 19573 9578 19625 9630
rect 19673 9060 19725 9112
rect 29701 8838 29753 8890
rect 29701 8468 29753 8520
rect 19573 8246 19625 8298
rect 19673 7728 19725 7780
rect 29701 7506 29753 7558
rect 29701 7136 29753 7188
rect 19573 6914 19625 6966
rect 10926 4116 13292 4314
rect 13684 3983 13736 4035
rect 10824 2034 13454 2234
rect 20254 1840 20306 1960
rect 20358 1840 20410 1960
rect 29086 1840 29138 1960
rect 29190 1840 29242 1960
<< metal2 >>
rect 20908 12377 20991 12386
rect 20908 12274 20991 12283
rect 20924 12158 20972 12274
rect 20649 12110 20972 12158
rect 19671 11704 19727 11714
rect 19671 11638 19727 11648
rect 29699 11556 29755 11566
rect 29699 11490 29755 11500
rect 29699 11186 29755 11196
rect 29699 11120 29755 11130
rect 19571 10964 19627 10974
rect 19571 10898 19627 10908
rect 19671 10446 19727 10456
rect 19671 10380 19727 10390
rect 29699 10224 29755 10234
rect 29699 10158 29755 10168
rect 29699 9854 29755 9864
rect 29699 9788 29755 9798
rect 19571 9632 19627 9642
rect 19571 9566 19627 9576
rect 19671 9114 19727 9124
rect 19671 9048 19727 9058
rect 29699 8892 29755 8902
rect 29699 8826 29755 8836
rect 29699 8522 29755 8532
rect 29699 8456 29755 8466
rect 19571 8300 19627 8310
rect 19571 8234 19627 8244
rect 19671 7782 19727 7792
rect 19671 7716 19727 7726
rect 29699 7560 29755 7570
rect 29699 7494 29755 7504
rect 29699 7190 29755 7200
rect 29699 7124 29755 7134
rect 19571 6968 19627 6978
rect 19571 6902 19627 6912
rect 19737 5200 23983 5248
rect 24345 5200 28617 5248
rect 19737 4592 19785 5200
rect 28569 4592 28617 5200
rect 10660 4488 10669 4571
rect 10763 4552 10772 4571
rect 10763 4504 10855 4552
rect 10763 4488 10772 4504
rect 10819 4374 10855 4504
rect 17688 4340 17958 4400
rect 26448 4340 26790 4400
rect 10920 4116 10926 4314
rect 13292 4116 13298 4314
rect 13684 4035 13736 4041
rect 13684 3965 13736 3983
rect 13667 3956 13750 3965
rect 13667 3853 13750 3862
rect 17688 2907 17740 4340
rect 13468 2855 17740 2907
rect 13468 2515 17740 2567
rect 10818 2034 10824 2234
rect 13454 2034 13460 2234
rect 17688 1572 17740 2515
rect 19994 1840 20003 1960
rect 20188 1840 20254 1960
rect 20306 1840 20312 1960
rect 20352 1840 20358 1960
rect 20410 1840 20476 1960
rect 20661 1840 20670 1960
rect 26448 1572 26500 4340
rect 28826 1840 28835 1960
rect 29020 1840 29086 1960
rect 29138 1840 29144 1960
rect 29184 1840 29190 1960
rect 29242 1840 29308 1960
rect 29493 1840 29502 1960
rect 17688 1520 26500 1572
<< via2 >>
rect 20908 12283 20991 12377
rect 19671 11702 19727 11704
rect 19671 11650 19673 11702
rect 19673 11650 19725 11702
rect 19725 11650 19727 11702
rect 19671 11648 19727 11650
rect 29699 11554 29755 11556
rect 29699 11502 29701 11554
rect 29701 11502 29753 11554
rect 29753 11502 29755 11554
rect 29699 11500 29755 11502
rect 29699 11184 29755 11186
rect 29699 11132 29701 11184
rect 29701 11132 29753 11184
rect 29753 11132 29755 11184
rect 29699 11130 29755 11132
rect 19571 10962 19627 10964
rect 19571 10910 19573 10962
rect 19573 10910 19625 10962
rect 19625 10910 19627 10962
rect 19571 10908 19627 10910
rect 19671 10444 19727 10446
rect 19671 10392 19673 10444
rect 19673 10392 19725 10444
rect 19725 10392 19727 10444
rect 19671 10390 19727 10392
rect 29699 10222 29755 10224
rect 29699 10170 29701 10222
rect 29701 10170 29753 10222
rect 29753 10170 29755 10222
rect 29699 10168 29755 10170
rect 29699 9852 29755 9854
rect 29699 9800 29701 9852
rect 29701 9800 29753 9852
rect 29753 9800 29755 9852
rect 29699 9798 29755 9800
rect 19571 9630 19627 9632
rect 19571 9578 19573 9630
rect 19573 9578 19625 9630
rect 19625 9578 19627 9630
rect 19571 9576 19627 9578
rect 19671 9112 19727 9114
rect 19671 9060 19673 9112
rect 19673 9060 19725 9112
rect 19725 9060 19727 9112
rect 19671 9058 19727 9060
rect 29699 8890 29755 8892
rect 29699 8838 29701 8890
rect 29701 8838 29753 8890
rect 29753 8838 29755 8890
rect 29699 8836 29755 8838
rect 29699 8520 29755 8522
rect 29699 8468 29701 8520
rect 29701 8468 29753 8520
rect 29753 8468 29755 8520
rect 29699 8466 29755 8468
rect 19571 8298 19627 8300
rect 19571 8246 19573 8298
rect 19573 8246 19625 8298
rect 19625 8246 19627 8298
rect 19571 8244 19627 8246
rect 19671 7780 19727 7782
rect 19671 7728 19673 7780
rect 19673 7728 19725 7780
rect 19725 7728 19727 7780
rect 19671 7726 19727 7728
rect 29699 7558 29755 7560
rect 29699 7506 29701 7558
rect 29701 7506 29753 7558
rect 29753 7506 29755 7558
rect 29699 7504 29755 7506
rect 29699 7188 29755 7190
rect 29699 7136 29701 7188
rect 29701 7136 29753 7188
rect 29753 7136 29755 7188
rect 29699 7134 29755 7136
rect 19571 6966 19627 6968
rect 19571 6914 19573 6966
rect 19573 6914 19625 6966
rect 19625 6914 19627 6966
rect 19571 6912 19627 6914
rect 10669 4488 10763 4571
rect 10929 4121 13289 4309
rect 13667 3862 13750 3956
rect 10827 2039 13451 2229
rect 20003 1840 20188 1960
rect 20476 1840 20661 1960
rect 28835 1840 29020 1960
rect 29308 1840 29493 1960
<< metal3 >>
rect 6682 44862 6750 44868
rect 6682 44798 6684 44862
rect 6748 44798 6750 44862
rect 6682 44792 6750 44798
rect 7418 44862 7486 44868
rect 7418 44798 7420 44862
rect 7484 44798 7486 44862
rect 7418 44792 7486 44798
rect 8154 44862 8222 44868
rect 8154 44798 8156 44862
rect 8220 44798 8222 44862
rect 8154 44792 8222 44798
rect 8890 44862 8958 44868
rect 8890 44798 8892 44862
rect 8956 44798 8958 44862
rect 8890 44792 8958 44798
rect 9626 44862 9694 44868
rect 9626 44798 9628 44862
rect 9692 44798 9694 44862
rect 9626 44792 9694 44798
rect 10362 44862 10430 44868
rect 10362 44798 10364 44862
rect 10428 44798 10430 44862
rect 10362 44792 10430 44798
rect 11098 44862 11166 44868
rect 11098 44798 11100 44862
rect 11164 44798 11166 44862
rect 11098 44792 11166 44798
rect 11834 44862 11902 44868
rect 11834 44798 11836 44862
rect 11900 44798 11902 44862
rect 11834 44792 11902 44798
rect 12570 44862 12638 44868
rect 12570 44798 12572 44862
rect 12636 44798 12638 44862
rect 12570 44792 12638 44798
rect 13306 44862 13374 44868
rect 13306 44798 13308 44862
rect 13372 44798 13374 44862
rect 13306 44792 13374 44798
rect 14042 44862 14110 44868
rect 14042 44798 14044 44862
rect 14108 44798 14110 44862
rect 14042 44792 14110 44798
rect 14778 44862 14846 44868
rect 14778 44798 14780 44862
rect 14844 44798 14846 44862
rect 14778 44792 14846 44798
rect 15514 44862 15582 44868
rect 15514 44798 15516 44862
rect 15580 44798 15582 44862
rect 15514 44792 15582 44798
rect 16250 44862 16318 44868
rect 16250 44798 16252 44862
rect 16316 44798 16318 44862
rect 16250 44792 16318 44798
rect 16986 44862 17054 44868
rect 16986 44798 16988 44862
rect 17052 44798 17054 44862
rect 16986 44792 17054 44798
rect 17722 44862 17790 44868
rect 17722 44798 17724 44862
rect 17788 44798 17790 44862
rect 17722 44792 17790 44798
rect 6686 42300 6746 44792
rect 7422 42460 7482 44792
rect 8158 42620 8218 44792
rect 8894 42780 8954 44792
rect 9630 42940 9690 44792
rect 10366 43100 10426 44792
rect 11102 43260 11162 44792
rect 11838 43420 11898 44792
rect 12574 43580 12634 44792
rect 13310 43740 13370 44792
rect 14046 43900 14106 44792
rect 14782 44060 14842 44792
rect 15518 44220 15578 44792
rect 16254 44380 16314 44792
rect 16990 44540 17050 44792
rect 17726 44700 17786 44792
rect 17726 44640 19567 44700
rect 16990 44480 19407 44540
rect 16254 44320 19247 44380
rect 15518 44160 19087 44220
rect 14782 44000 18927 44060
rect 14046 43840 18767 43900
rect 13310 43680 18607 43740
rect 12574 43520 18447 43580
rect 11838 43360 18287 43420
rect 11102 43200 18127 43260
rect 10366 43040 17967 43100
rect 9630 42880 17807 42940
rect 8894 42720 17647 42780
rect 8158 42560 17487 42620
rect 7422 42400 17327 42460
rect 6686 42240 17167 42300
rect 17107 6810 17167 42240
rect 17267 6970 17327 42400
rect 17427 7562 17487 42560
rect 17587 7784 17647 42720
rect 17747 8142 17807 42880
rect 17907 8302 17967 43040
rect 18067 8894 18127 43200
rect 18227 9116 18287 43360
rect 18387 9474 18447 43520
rect 18547 9634 18607 43680
rect 18707 10226 18767 43840
rect 18867 10448 18927 44000
rect 19027 10806 19087 44160
rect 19187 10966 19247 44320
rect 19347 11558 19407 44480
rect 19507 11706 19567 44640
rect 20902 12377 20997 12383
rect 20902 12283 20908 12377
rect 20991 12283 20997 12377
rect 20902 12277 20997 12283
rect 19665 11706 19733 11710
rect 19507 11704 19733 11706
rect 19507 11648 19671 11704
rect 19727 11648 19733 11704
rect 19507 11646 19733 11648
rect 19665 11642 19733 11646
rect 29693 11558 29761 11562
rect 19347 11556 29761 11558
rect 19347 11500 29699 11556
rect 29755 11500 29761 11556
rect 19347 11498 29761 11500
rect 29693 11494 29761 11498
rect 29693 11188 29761 11192
rect 19713 11186 29761 11188
rect 19713 11130 29699 11186
rect 29755 11130 29761 11186
rect 19713 11128 29761 11130
rect 19565 10966 19633 10970
rect 19187 10964 19633 10966
rect 19187 10908 19571 10964
rect 19627 10908 19633 10964
rect 19187 10906 19633 10908
rect 19565 10902 19633 10906
rect 19713 10806 19773 11128
rect 29693 11124 29761 11128
rect 19027 10746 19773 10806
rect 19665 10448 19733 10452
rect 18867 10446 19733 10448
rect 18867 10390 19671 10446
rect 19727 10390 19733 10446
rect 18867 10388 19733 10390
rect 19665 10384 19733 10388
rect 29693 10226 29761 10230
rect 18707 10224 29761 10226
rect 18707 10168 29699 10224
rect 29755 10168 29761 10224
rect 18707 10166 29761 10168
rect 29693 10162 29761 10166
rect 29693 9856 29761 9860
rect 19713 9854 29761 9856
rect 19713 9798 29699 9854
rect 29755 9798 29761 9854
rect 19713 9796 29761 9798
rect 19565 9634 19633 9638
rect 18547 9632 19633 9634
rect 18547 9576 19571 9632
rect 19627 9576 19633 9632
rect 18547 9574 19633 9576
rect 19565 9570 19633 9574
rect 19713 9474 19773 9796
rect 29693 9792 29761 9796
rect 18387 9414 19773 9474
rect 19665 9116 19733 9120
rect 18227 9114 19733 9116
rect 18227 9058 19671 9114
rect 19727 9058 19733 9114
rect 18227 9056 19733 9058
rect 19665 9052 19733 9056
rect 29693 8894 29761 8898
rect 18067 8892 29761 8894
rect 18067 8836 29699 8892
rect 29755 8836 29761 8892
rect 18067 8834 29761 8836
rect 29693 8830 29761 8834
rect 29693 8524 29761 8528
rect 19713 8522 29761 8524
rect 19713 8466 29699 8522
rect 29755 8466 29761 8522
rect 19713 8464 29761 8466
rect 19565 8302 19633 8306
rect 17907 8300 19633 8302
rect 17907 8244 19571 8300
rect 19627 8244 19633 8300
rect 17907 8242 19633 8244
rect 19565 8238 19633 8242
rect 19713 8142 19773 8464
rect 29693 8460 29761 8464
rect 17747 8082 19773 8142
rect 19665 7784 19733 7788
rect 17587 7782 19733 7784
rect 17587 7726 19671 7782
rect 19727 7726 19733 7782
rect 17587 7724 19733 7726
rect 19665 7720 19733 7724
rect 29693 7562 29761 7566
rect 17427 7560 29761 7562
rect 17427 7504 29699 7560
rect 29755 7504 29761 7560
rect 17427 7502 29761 7504
rect 29693 7498 29761 7502
rect 29693 7192 29761 7196
rect 19713 7190 29761 7192
rect 19713 7134 29699 7190
rect 29755 7134 29761 7190
rect 19713 7132 29761 7134
rect 19565 6970 19633 6974
rect 17267 6968 19633 6970
rect 17267 6912 19571 6968
rect 19627 6912 19633 6968
rect 17267 6910 19633 6912
rect 19565 6906 19633 6910
rect 19713 6810 19773 7132
rect 29693 7128 29761 7132
rect 17107 6750 19773 6810
rect 10663 4571 10769 4577
rect 10663 4488 10669 4571
rect 10763 4488 10769 4571
rect 10663 4482 10769 4488
rect 10920 4313 13298 4314
rect 10920 4309 12061 4313
rect 12359 4309 13298 4313
rect 10920 4121 10929 4309
rect 13289 4121 13298 4309
rect 10920 4117 12061 4121
rect 12359 4117 13298 4121
rect 10920 4116 13298 4117
rect 13661 3956 13756 3962
rect 13661 3862 13667 3956
rect 13750 3862 13756 3956
rect 13661 3856 13756 3862
rect 20205 2579 20550 2580
rect 10818 2233 13460 2234
rect 10818 2229 11661 2233
rect 11959 2229 13460 2233
rect 10818 2039 10827 2229
rect 13451 2039 13460 2229
rect 20205 2081 20306 2579
rect 20544 2081 20550 2579
rect 20205 2080 20550 2081
rect 29037 2579 29509 2580
rect 29037 2081 29265 2579
rect 29503 2081 29509 2579
rect 29037 2080 29509 2081
rect 10818 2035 11661 2039
rect 11959 2035 13460 2039
rect 10818 2034 13460 2035
rect 19998 1960 20193 1965
rect 18064 1840 20003 1960
rect 20188 1840 20193 1960
rect 18064 394 18184 1840
rect 19998 1835 20193 1840
rect 20471 1960 20666 1965
rect 28830 1960 29025 1965
rect 20471 1840 20476 1960
rect 20661 1840 22600 1960
rect 20471 1835 20666 1840
rect 18064 200 18184 206
rect 22480 394 22600 1840
rect 22480 200 22600 206
rect 26896 1840 28835 1960
rect 29020 1840 29025 1960
rect 26896 394 27016 1840
rect 28830 1835 29025 1840
rect 29303 1960 29498 1965
rect 29303 1840 29308 1960
rect 29493 1840 31432 1960
rect 29303 1835 29498 1840
rect 26896 200 27016 206
rect 31312 394 31432 1840
rect 31312 200 31432 206
<< via3 >>
rect 6684 44798 6748 44862
rect 7420 44798 7484 44862
rect 8156 44798 8220 44862
rect 8892 44798 8956 44862
rect 9628 44798 9692 44862
rect 10364 44798 10428 44862
rect 11100 44798 11164 44862
rect 11836 44798 11900 44862
rect 12572 44798 12636 44862
rect 13308 44798 13372 44862
rect 14044 44798 14108 44862
rect 14780 44798 14844 44862
rect 15516 44798 15580 44862
rect 16252 44798 16316 44862
rect 16988 44798 17052 44862
rect 17724 44798 17788 44862
rect 20918 12298 20982 12362
rect 10684 4498 10748 4562
rect 12061 4309 12359 4313
rect 12061 4121 12359 4309
rect 12061 4117 12359 4121
rect 13676 3877 13740 3941
rect 18561 3377 19999 3503
rect 27393 3377 28831 3503
rect 11661 2229 11959 2233
rect 11661 2039 11959 2229
rect 20306 2081 20544 2579
rect 29265 2081 29503 2579
rect 11661 2035 11959 2039
rect 18064 206 18184 394
rect 22480 206 22600 394
rect 26896 206 27016 394
rect 31312 206 31432 394
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 440 44892 6010 44952
rect 440 44152 500 44892
rect 6686 44864 6746 45152
rect 7422 44864 7482 45152
rect 8158 44864 8218 45152
rect 8894 44864 8954 45152
rect 9630 44864 9690 45152
rect 10366 44864 10426 45152
rect 11102 44864 11162 45152
rect 11838 44864 11898 45152
rect 12574 44864 12634 45152
rect 13310 44864 13370 45152
rect 14046 44864 14106 45152
rect 14782 44864 14842 45152
rect 15518 44864 15578 45152
rect 16254 44864 16314 45152
rect 16990 44864 17050 45152
rect 17726 44864 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 6682 44862 6750 44864
rect 6682 44798 6684 44862
rect 6748 44798 6750 44862
rect 6682 44796 6750 44798
rect 7418 44862 7486 44864
rect 7418 44798 7420 44862
rect 7484 44798 7486 44862
rect 7418 44796 7486 44798
rect 8154 44862 8222 44864
rect 8154 44798 8156 44862
rect 8220 44798 8222 44862
rect 8154 44796 8222 44798
rect 8890 44862 8958 44864
rect 8890 44798 8892 44862
rect 8956 44798 8958 44862
rect 8890 44796 8958 44798
rect 9626 44862 9694 44864
rect 9626 44798 9628 44862
rect 9692 44798 9694 44862
rect 9626 44796 9694 44798
rect 10362 44862 10430 44864
rect 10362 44798 10364 44862
rect 10428 44798 10430 44862
rect 10362 44796 10430 44798
rect 11098 44862 11166 44864
rect 11098 44798 11100 44862
rect 11164 44798 11166 44862
rect 11098 44796 11166 44798
rect 11834 44862 11902 44864
rect 11834 44798 11836 44862
rect 11900 44798 11902 44862
rect 11834 44796 11902 44798
rect 12570 44862 12638 44864
rect 12570 44798 12572 44862
rect 12636 44798 12638 44862
rect 12570 44796 12638 44798
rect 13306 44862 13374 44864
rect 13306 44798 13308 44862
rect 13372 44798 13374 44862
rect 13306 44796 13374 44798
rect 14042 44862 14110 44864
rect 14042 44798 14044 44862
rect 14108 44798 14110 44862
rect 14042 44796 14110 44798
rect 14778 44862 14846 44864
rect 14778 44798 14780 44862
rect 14844 44798 14846 44862
rect 14778 44796 14846 44798
rect 15514 44862 15582 44864
rect 15514 44798 15516 44862
rect 15580 44798 15582 44862
rect 15514 44796 15582 44798
rect 16250 44862 16318 44864
rect 16250 44798 16252 44862
rect 16316 44798 16318 44862
rect 16250 44796 16318 44798
rect 16986 44862 17054 44864
rect 16986 44798 16988 44862
rect 17052 44798 17054 44862
rect 16986 44796 17054 44798
rect 17722 44862 17790 44864
rect 17722 44798 17724 44862
rect 17788 44798 17790 44862
rect 17722 44796 17790 44798
rect 28766 44420 28826 45152
rect 9460 44360 28826 44420
rect 8040 44152 8100 44200
rect 200 1000 500 44152
rect 600 23300 900 44152
rect 7800 29100 8100 44152
rect 600 22900 1500 23300
rect 600 17000 900 22900
rect 600 16600 1500 17000
rect 600 10600 900 16600
rect 600 10200 1500 10600
rect 600 1000 900 10200
rect 7700 10000 8100 29100
rect 7800 1000 8100 10000
rect 9460 4560 9520 44360
rect 29502 44280 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 20920 44220 29562 44280
rect 10683 4562 10749 4563
rect 10683 4560 10684 4562
rect 9460 4500 10684 4560
rect 10683 4498 10684 4500
rect 10748 4498 10749 4562
rect 10683 4497 10749 4498
rect 11660 2233 11960 44152
rect 11660 2035 11661 2233
rect 11959 2035 11960 2233
rect 11660 1000 11960 2035
rect 12060 4313 12360 44152
rect 12060 4117 12061 4313
rect 12359 4117 12360 4313
rect 12060 1000 12360 4117
rect 13675 3941 13741 3942
rect 13675 3877 13676 3941
rect 13740 3877 13741 3941
rect 13675 3840 13741 3877
rect 13648 200 13768 3840
rect 19845 3504 20145 44152
rect 18555 3503 20145 3504
rect 18555 3377 18561 3503
rect 19999 3377 20145 3503
rect 18555 3376 20145 3377
rect 19845 1000 20145 3376
rect 20305 2579 20605 44152
rect 20920 12363 20980 44220
rect 20917 12362 20983 12363
rect 20917 12298 20918 12362
rect 20982 12298 20983 12362
rect 20917 12297 20983 12298
rect 28804 3504 29104 44152
rect 27387 3503 29104 3504
rect 27387 3377 27393 3503
rect 28831 3377 29104 3503
rect 27387 3376 29104 3377
rect 20305 2081 20306 2579
rect 20544 2081 20605 2579
rect 20305 1000 20605 2081
rect 28804 1000 29104 3376
rect 29264 2579 29564 44152
rect 29264 2081 29265 2579
rect 29503 2081 29564 2579
rect 29264 1000 29564 2081
rect 18034 394 18214 400
rect 18034 206 18064 394
rect 18184 206 18214 394
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 206
rect 22450 394 22630 400
rect 22450 206 22480 394
rect 22600 206 22630 394
rect 22450 0 22630 206
rect 26866 394 27046 400
rect 26866 206 26896 394
rect 27016 206 27046 394
rect 26866 0 27046 206
rect 31282 394 31462 400
rect 31282 206 31312 394
rect 31432 206 31462 394
rect 31282 0 31462 206
use bias_gen  bias_gen_0 usb
timestamp 1717081332
transform 0 1 10360 -1 0 5154
box 780 -360 3154 3160
use diff_rx  diff_rx_0 usb
timestamp 1717246753
transform 1 0 18618 0 1 2100
box -720 -100 3488 2767
use diff_rx  diff_rx_1
timestamp 1717246753
transform 1 0 27450 0 1 2100
box -720 -100 3488 2767
use digital  digital_0 usb
timestamp 1717248114
transform 1 0 25761 0 1 7347
box -5994 -2147 3898 4811
use sky130_fd_pr__cap_mim_m3_1_L66JLG  sky130_fd_pr__cap_mim_m3_1_L66JLG_0
timestamp 1717266104
transform 1 0 4586 0 1 19480
box -3186 -9480 3186 9480
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 5 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 53 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 52 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 51 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 50 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 49 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 48 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 47 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 46 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 13 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 11 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 10 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 7 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 6 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 21 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 19 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 18 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 15 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 14 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 45 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 44 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 43 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 42 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 41 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 40 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 39 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 37 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 35 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 34 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 31 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 30 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 29 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 28 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 27 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 26 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 25 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 24 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 23 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 22 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 720 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 600 1000 900 44152 1 FreeSans 720 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 38 nsew signal output
flabel metal4 19845 1000 20145 44152 0 FreeSans 320 0 0 0 VGND
port 1 nsew
flabel metal4 20305 1000 20605 44152 0 FreeSans 320 0 0 0 VPWR
port 2 nsew
flabel metal4 28804 1000 29104 44152 0 FreeSans 320 0 0 0 VGND
port 1 nsew
flabel metal4 29264 1000 29564 44152 0 FreeSans 320 0 0 0 VPWR
port 2 nsew
flabel metal4 11660 1000 11960 44152 1 FreeSans 720 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 12060 1000 12360 44152 1 FreeSans 720 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 7800 1000 8100 44152 1 FreeSans 720 0 0 0 VPWR
port 2 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
